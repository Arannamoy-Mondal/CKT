CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 880 30 100 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 138 1416 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3835 0 0
2
45780 0
0
13 Logic Switch~
5 138 1334 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3670 0 0
2
45780 0
0
13 Logic Switch~
5 135 1256 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5616 0 0
2
45780 0
0
13 Logic Switch~
5 172 349 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9323 0 0
2
45779.9 0
0
13 Logic Switch~
5 169 282 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
317 0 0
2
45779.9 0
0
13 Logic Switch~
5 172 206 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3108 0 0
2
45779.9 0
0
9 Inverter~
13 215 1375 0 2 22
0 7 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
4299 0 0
2
45780 0
0
14 Logic Display~
6 653 1323 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9672 0 0
2
45780 0
0
5 4071~
219 478 1329 0 3 22
0 4 3 2
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
7876 0 0
2
45780 0
0
5 4081~
219 335 1393 0 3 22
0 6 5 3
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
6369 0 0
2
45780 0
0
5 4081~
219 331 1286 0 3 22
0 7 8 4
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
9172 0 0
2
45780 0
0
14 Logic Display~
6 749 520 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7100 0 0
2
45779.9 0
0
5 4071~
219 602 524 0 3 22
0 11 10 9
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
3820 0 0
2
45779.9 0
0
5 4081~
219 359 560 0 3 22
0 13 12 10
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
7678 0 0
2
45779.9 0
0
5 4081~
219 408 469 0 3 22
0 15 14 11
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
961 0 0
2
45779.9 0
0
14 Logic Display~
6 606 337 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3178 0 0
2
45779.9 0
0
9 2-In XOR~
219 415 339 0 3 22
0 15 14 16
0
0 0 624 0
7 74LS386
-24 -24 25 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3409 0 0
2
45779.9 0
0
9 2-In XOR~
219 331 233 0 3 22
0 13 12 15
0
0 0 624 0
7 74LS386
-24 -24 25 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3951 0 0
2
45779.9 0
0
20
3 1 2 0 0 4224 0 9 8 0 0 5
511 1329
641 1329
641 1349
653 1349
653 1341
3 2 3 0 0 4224 0 10 9 0 0 4
356 1393
457 1393
457 1338
465 1338
3 1 4 0 0 4224 0 11 9 0 0 4
352 1286
457 1286
457 1320
465 1320
1 2 5 0 0 4224 0 1 10 0 0 4
150 1416
303 1416
303 1402
311 1402
2 1 6 0 0 4224 0 7 10 0 0 4
236 1375
303 1375
303 1384
311 1384
0 1 7 0 0 4096 0 0 7 8 0 3
171 1256
171 1375
200 1375
1 2 8 0 0 4224 0 2 11 0 0 4
150 1334
299 1334
299 1295
307 1295
1 1 7 0 0 4224 0 3 11 0 0 4
147 1256
299 1256
299 1277
307 1277
3 1 9 0 0 4224 0 13 12 0 0 5
635 524
737 524
737 546
749 546
749 538
3 2 10 0 0 4224 0 14 13 0 0 4
380 560
581 560
581 533
589 533
3 1 11 0 0 4224 0 15 13 0 0 4
429 469
581 469
581 515
589 515
0 2 12 0 0 4224 0 0 14 19 0 3
196 282
196 569
335 569
0 1 13 0 0 4224 0 0 14 20 0 3
268 206
268 551
335 551
0 2 14 0 0 8192 0 0 15 17 0 3
251 349
251 478
384 478
0 1 15 0 0 4224 0 0 15 18 0 3
372 233
372 460
384 460
3 1 16 0 0 4224 0 17 16 0 0 5
448 339
594 339
594 363
606 363
606 355
1 2 14 0 0 4224 0 4 17 0 0 4
184 349
391 349
391 348
399 348
3 1 15 0 0 128 0 18 17 0 0 4
364 233
391 233
391 330
399 330
1 2 12 0 0 128 0 5 18 0 0 4
181 282
307 282
307 242
315 242
1 1 13 0 0 128 0 6 18 0 0 4
184 206
307 206
307 224
315 224
13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
50 1400 87 1424
60 1408 76 1424
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
54 1326 91 1350
64 1334 80 1350
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
52 1237 89 1261
62 1245 78 1261
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
63 1095 116 1119
73 1103 105 1119
4 2.b)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
632 485 741 509
642 493 730 509
11 C(A(+)B)+AB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
401 526 438 550
411 534 427 550
2 AB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
432 429 517 453
442 437 506 453
8 c(A(+)B)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
464 298 557 322
474 306 546 322
9 A(+)B(+)C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
360 178 421 202
370 186 410 202
5 A(+)B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
102 325 127 349
110 333 118 349
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
109 263 138 287
119 271 127 287
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
127 186 156 210
137 194 145 210
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
74 48 127 72
84 56 116 72
4 2.a)
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
