CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 1180 30 100 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
49
13 Logic Switch~
5 108 1683 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V21
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4299 0 0
2
45780.1 0
0
13 Logic Switch~
5 108 1638 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V20
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9672 0 0
2
45780.1 0
0
13 Logic Switch~
5 109 1593 0 1 11
0 7
0
0 0 21360 0
2 0V
-4 -15 10 -7
3 V19
-8 -24 13 -16
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7876 0 0
2
45780.1 0
0
13 Logic Switch~
5 108 1558 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V18
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6369 0 0
2
45780.1 0
0
13 Logic Switch~
5 109 1524 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V17
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9172 0 0
2
45780.1 0
0
13 Logic Switch~
5 112 1487 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V16
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7100 0 0
2
45780.1 0
0
13 Logic Switch~
5 105 1453 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V15
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3820 0 0
2
45780.1 0
0
13 Logic Switch~
5 106 1412 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V14
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7678 0 0
2
45780.1 0
0
13 Logic Switch~
5 104 1371 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V13
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
961 0 0
2
45780.1 0
0
13 Logic Switch~
5 80 1108 0 1 11
0 25
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3178 0 0
2
45780.1 0
0
13 Logic Switch~
5 73 1079 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3409 0 0
2
45780.1 0
0
13 Logic Switch~
5 72 1037 0 1 11
0 27
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3951 0 0
2
45780.1 0
0
13 Logic Switch~
5 69 995 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8885 0 0
2
45780.1 0
0
13 Logic Switch~
5 60 951 0 1 11
0 29
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3780 0 0
2
45780.1 0
0
13 Logic Switch~
5 59 908 0 10 11
0 30 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9265 0 0
2
45780.1 0
0
13 Logic Switch~
5 57 869 0 1 11
0 31
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9442 0 0
2
45780.1 0
0
13 Logic Switch~
5 61 823 0 10 11
0 32 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9424 0 0
2
45780.1 0
0
13 Logic Switch~
5 65 776 0 10 11
0 33 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-5 -27 9 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9968 0 0
2
45780.1 0
0
13 Logic Switch~
5 86 321 0 10 11
0 39 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9281 0 0
2
45780 0
0
13 Logic Switch~
5 87 179 0 10 11
0 41 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8464 0 0
2
45780 0
0
13 Logic Switch~
5 90 121 0 10 11
0 40 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7168 0 0
2
45780 0
0
9 Inverter~
13 170 1636 0 2 22
0 6 2
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 5 0
1 U
3171 0 0
2
45780.1 0
0
9 Inverter~
13 172 1591 0 2 22
0 7 3
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 5 0
1 U
4139 0 0
2
45780.1 0
0
9 Inverter~
13 173 1557 0 2 22
0 8 4
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 5 0
1 U
6435 0 0
2
45780.1 0
0
9 Inverter~
13 172 1526 0 2 22
0 9 5
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 5 0
1 U
5283 0 0
2
45780.1 0
0
14 Logic Display~
6 502 1604 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L14
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6874 0 0
2
45780.1 0
0
14 Logic Display~
6 504 1550 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5305 0 0
2
45780.1 0
0
14 Logic Display~
6 501 1491 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
34 0 0
2
45780.1 0
0
14 Logic Display~
6 501 1435 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
969 0 0
2
45780.1 0
0
14 Logic Display~
6 500 1372 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8402 0 0
2
45780.1 0
0
6 74LS83
105 303 1419 0 14 29
0 18 19 10 11 2 3 4 5 17
13 14 15 16 12
0
0 0 4848 0
7 74LS83A
-24 -60 25 -52
2 U6
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 0 0 0 0
1 U
3751 0 0
2
45780.1 0
0
14 Logic Display~
6 496 1007 0 1 2
10 20
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4292 0 0
2
45780.1 0
0
14 Logic Display~
6 493 962 0 1 2
10 21
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6118 0 0
2
45780.1 0
0
14 Logic Display~
6 489 917 0 1 2
10 22
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
34 0 0
2
45780.1 0
0
14 Logic Display~
6 489 867 0 1 2
10 23
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6357 0 0
2
45780.1 0
0
14 Logic Display~
6 487 821 0 1 2
10 24
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
319 0 0
2
45780.1 0
0
6 74LS83
105 280 850 0 14 29
0 30 31 32 33 26 27 28 29 25
21 22 23 24 20
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U5
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 0 0 0 0
1 U
3976 0 0
2
45780.1 0
0
5 4071~
219 374 441 0 3 22
0 36 35 34
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
7634 0 0
2
45780.1 0
0
5 4071~
219 286 427 0 3 22
0 38 37 36
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
523 0 0
2
45780.1 0
0
5 4081~
219 202 545 0 3 22
0 40 39 35
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
6748 0 0
2
45780.1 0
0
5 4081~
219 214 468 0 3 22
0 41 39 37
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
6901 0 0
2
45780.1 0
0
5 4081~
219 203 400 0 3 22
0 40 41 38
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
842 0 0
2
45780.1 0
0
14 Logic Display~
6 434 392 0 1 2
10 34
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3277 0 0
2
45780.1 0
0
14 Logic Display~
6 432 319 0 1 2
10 42
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4212 0 0
2
45780.1 0
0
9 2-In XOR~
219 297 313 0 3 22
0 43 39 42
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U3A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
4720 0 0
2
45780 0
0
14 Logic Display~
6 386 213 0 1 2
10 44
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5551 0 0
2
45780 0
0
14 Logic Display~
6 383 139 0 1 2
10 43
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6986 0 0
2
45780 0
0
5 4081~
219 208 220 0 3 22
0 40 41 44
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
8745 0 0
2
45780 0
0
9 2-In XOR~
219 216 137 0 3 22
0 40 41 43
0
0 0 624 0
7 74LS386
-24 -24 25 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9592 0 0
2
45780 0
0
52
2 5 2 0 0 8320 0 22 31 0 0 4
191 1636
238 1636
238 1419
271 1419
2 6 3 0 0 8320 0 23 31 0 0 4
193 1591
243 1591
243 1428
271 1428
2 7 4 0 0 8336 0 24 31 0 0 4
194 1557
258 1557
258 1437
271 1437
2 8 5 0 0 8320 0 25 31 0 0 4
193 1526
263 1526
263 1446
271 1446
1 1 6 0 0 4224 0 2 22 0 0 4
120 1638
147 1638
147 1636
155 1636
1 1 7 0 0 4224 0 3 23 0 0 4
121 1593
149 1593
149 1591
157 1591
1 1 8 0 0 4224 0 4 24 0 0 4
120 1558
150 1558
150 1557
158 1557
1 1 9 0 0 4224 0 5 25 0 0 4
121 1524
149 1524
149 1526
157 1526
1 3 10 0 0 4224 0 8 31 0 0 4
118 1412
258 1412
258 1401
271 1401
1 4 11 0 0 4224 0 9 31 0 0 4
116 1371
263 1371
263 1410
271 1410
14 1 12 0 0 4224 0 31 26 0 0 8
335 1464
335 1627
439 1627
439 1625
484 1625
484 1630
502 1630
502 1622
10 1 13 0 0 8320 0 31 27 0 0 7
335 1410
421 1410
421 1535
491 1535
491 1576
504 1576
504 1568
11 1 14 0 0 4224 0 31 28 0 0 5
335 1419
478 1419
478 1517
501 1517
501 1509
12 1 15 0 0 4224 0 31 29 0 0 5
335 1428
484 1428
484 1461
501 1461
501 1453
13 1 16 0 0 4224 0 31 30 0 0 5
335 1437
489 1437
489 1398
500 1398
500 1390
1 9 17 0 0 8320 0 1 31 0 0 4
120 1683
253 1683
253 1464
271 1464
1 1 18 0 0 4224 0 6 31 0 0 4
124 1487
248 1487
248 1383
271 1383
1 2 19 0 0 4224 0 7 31 0 0 4
117 1453
253 1453
253 1392
271 1392
14 1 20 0 0 8320 0 37 32 0 0 6
312 895
312 1071
586 1071
586 1022
496 1022
496 1025
10 1 21 0 0 4224 0 37 33 0 0 5
312 841
460 841
460 988
493 988
493 980
11 1 22 0 0 4224 0 37 34 0 0 5
312 850
466 850
466 943
489 943
489 935
12 1 23 0 0 4224 0 37 35 0 0 5
312 859
472 859
472 893
489 893
489 885
13 1 24 0 0 8320 0 37 36 0 0 6
312 868
312 825
477 825
477 847
487 847
487 839
1 9 25 0 0 8320 0 10 37 0 0 4
92 1108
226 1108
226 895
248 895
1 5 26 0 0 8320 0 11 37 0 0 4
85 1079
211 1079
211 850
248 850
1 6 27 0 0 8320 0 12 37 0 0 4
84 1037
216 1037
216 859
248 859
1 7 28 0 0 4224 0 13 37 0 0 4
81 995
231 995
231 868
248 868
1 8 29 0 0 4224 0 14 37 0 0 4
72 951
236 951
236 877
248 877
1 1 30 0 0 4224 0 15 37 0 0 4
71 908
221 908
221 814
248 814
1 2 31 0 0 4224 0 16 37 0 0 4
69 869
226 869
226 823
248 823
1 3 32 0 0 4224 0 17 37 0 0 4
73 823
231 823
231 832
248 832
1 4 33 0 0 4224 0 18 37 0 0 4
77 776
236 776
236 841
248 841
3 1 34 0 0 8320 0 38 43 0 0 3
407 441
434 441
434 410
3 2 35 0 0 4224 0 40 38 0 0 4
223 545
353 545
353 450
361 450
3 1 36 0 0 4224 0 39 38 0 0 4
319 427
353 427
353 432
361 432
3 2 37 0 0 8320 0 41 39 0 0 4
235 468
265 468
265 436
273 436
3 1 38 0 0 4224 0 42 39 0 0 4
224 400
265 400
265 418
273 418
0 2 39 0 0 4096 0 0 40 40 0 5
174 477
174 526
170 526
170 554
178 554
0 1 40 0 0 4096 0 0 40 43 0 3
158 391
158 536
178 536
0 2 39 0 0 4096 0 0 41 45 0 3
174 321
174 477
190 477
0 1 41 0 0 8192 0 0 41 42 0 3
132 409
132 459
190 459
0 2 41 0 0 4224 0 0 42 51 0 3
112 179
112 409
179 409
0 1 40 0 0 4224 0 0 42 52 0 3
143 121
143 391
179 391
3 1 42 0 0 4224 0 45 44 0 0 5
330 313
420 313
420 345
432 345
432 337
1 2 39 0 0 4224 0 19 45 0 0 4
98 321
273 321
273 322
281 322
0 1 43 0 0 4224 0 0 45 50 0 3
273 137
273 304
281 304
3 1 44 0 0 4224 0 48 46 0 0 5
229 220
374 220
374 239
386 239
386 231
0 2 41 0 0 0 0 0 48 51 0 3
158 179
158 229
184 229
0 1 40 0 0 128 0 0 48 52 0 3
128 121
128 211
184 211
3 1 43 0 0 128 0 49 47 0 0 5
249 137
371 137
371 165
383 165
383 157
1 2 41 0 0 128 0 20 49 0 0 4
99 179
192 179
192 146
200 146
1 1 40 0 0 128 0 21 49 0 0 4
102 121
192 121
192 128
200 128
40
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
39 1618 76 1642
49 1626 65 1642
2 B4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
53 1584 90 1608
63 1592 79 1608
2 B3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
48 1549 85 1573
58 1557 74 1573
2 B2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
39 1514 76 1538
49 1522 65 1538
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
31 1475 68 1499
41 1483 57 1499
2 A4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
16 1435 53 1459
26 1443 42 1459
2 A3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
22 1403 59 1427
32 1411 48 1427
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
18 1359 55 1383
28 1367 44 1383
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
48 1682 85 1706
58 1690 74 1706
2 Ci
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
545 1595 582 1619
555 1603 571 1619
2 Co
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
542 1538 579 1562
552 1546 568 1562
2 S4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
531 1477 568 1501
541 1485 557 1501
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
539 1425 576 1449
549 1433 565 1449
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
527 1363 564 1387
537 1371 553 1387
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 28
23 1216 268 1240
33 1224 257 1240
28 4.c)4 bit parallel Subtrator
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
25 1099 62 1123
35 1107 51 1123
2 Ci
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
534 987 571 1011
544 995 560 1011
2 C0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
527 943 564 967
537 951 553 967
2 S4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
516 901 553 925
526 909 542 925
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
528 850 565 874
538 858 554 874
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
513 802 550 826
523 810 539 826
2 s1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
5 1067 42 1091
15 1075 31 1091
2 B4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
11 1028 48 1052
21 1036 37 1052
2 B3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
13 988 50 1012
23 996 39 1012
2 B2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
9 930 46 954
19 938 35 954
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
11 888 48 912
21 896 37 912
2 A4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
10 841 47 865
20 849 36 865
2 A3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
15 799 52 823
25 807 41 823
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
9 764 46 788
19 772 35 788
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 24
30 690 243 714
40 698 232 714
24 4.b)4 bit Parallel Adder
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
331 371 432 395
341 379 421 395
10 C=AB+BC+AC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
511 307 628 331
521 315 617 331
12 (Full Adder)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
324 272 433 296
334 280 422 296
11 S=A(+)B(+)C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
21 297 50 321
31 305 39 321
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
217 178 270 202
227 186 259 202
4 C=AB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
432 119 549 143
442 127 538 143
12 (Half Adder)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
251 76 328 100
261 84 317 100
7 S=A(+)B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
28 146 57 170
38 154 46 170
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
29 85 58 109
39 93 47 109
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 40
24 0 229 44
34 8 218 40
40 4.a)Design Half Adder & 
    Full Adder
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
