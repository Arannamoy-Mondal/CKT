CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 1910 2 100 10
176 80 1278 731
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
57
13 Logic Switch~
5 190 1780 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V19
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3679 0 0
2
45781 2
0
13 Logic Switch~
5 179 1837 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V18
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9342 0 0
2
45781 1
0
13 Logic Switch~
5 175 1881 0 1 11
0 45
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V17
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 0 0 -2 0
1 V
3623 0 0
2
45781 0
0
13 Logic Switch~
5 140 1513 0 1 11
0 46
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V15
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 0 0 -2 0
1 V
3722 0 0
2
45781 2
0
13 Logic Switch~
5 144 1469 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V14
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8993 0 0
2
45781 1
0
13 Logic Switch~
5 155 1412 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V13
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3723 0 0
2
45781 0
0
13 Logic Switch~
5 192 1063 0 1 11
0 47
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V11
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 0 0 -2 0
1 V
6244 0 0
2
45781 2
0
13 Logic Switch~
5 196 1019 0 10 11
0 29 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6421 0 0
2
45781 1
0
13 Logic Switch~
5 207 962 0 10 11
0 30 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7743 0 0
2
45781 0
0
13 Logic Switch~
5 167 505 0 10 11
0 37 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9840 0 0
2
45781 2
0
13 Logic Switch~
5 156 562 0 10 11
0 36 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6910 0 0
2
45781 1
0
13 Logic Switch~
5 152 606 0 1 11
0 48
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 0 0 -2 0
1 V
449 0 0
2
45781 0
0
13 Logic Switch~
5 98 217 0 1 11
0 49
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 0 0 -2 0
1 V
8761 0 0
2
45781 0
0
13 Logic Switch~
5 102 173 0 10 11
0 43 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6748 0 0
2
45781 0
0
13 Logic Switch~
5 113 116 0 10 11
0 44 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7393 0 0
2
45781 0
0
5 4011~
219 876 1723 0 3 22
0 4 3 2
0
0 0 624 180
4 4011
-7 -24 21 -16
3 U5C
-8 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 5 0
1 U
7699 0 0
2
45781 0
0
14 Logic Display~
6 943 1986 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L16
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6638 0 0
2
45781 0
0
6 74112~
219 852 1827 0 7 32
0 2 8 5 8 7 3 6
0
0 0 4720 0
5 74112
4 -60 39 -52
4 U10B
19 -61 47 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 2 10 0
1 U
4595 0 0
2
45781 0
0
6 74112~
219 360 1833 0 7 32
0 2 8 13 8 7 12 11
0
0 0 4720 0
5 74112
4 -60 39 -52
4 U10A
19 -61 47 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 10 0
1 U
9395 0 0
2
45781 10
0
6 74112~
219 524 1827 0 7 32
0 2 8 12 8 7 4 10
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U9B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 2 9 0
1 U
3303 0 0
2
45781 9
0
6 74112~
219 677 1824 0 7 32
0 2 8 4 8 7 5 9
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U9A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 9 0
1 U
4498 0 0
2
45781 8
0
14 Logic Display~
6 450 2001 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L15
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9728 0 0
2
45781 7
0
14 Logic Display~
6 612 1995 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3789 0 0
2
45781 6
0
14 Logic Display~
6 801 1975 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3978 0 0
2
45781 5
0
7 Pulser~
4 172 2013 0 10 12
0 50 51 52 13 0 0 5 5 6
7
0
0 0 4656 0
0
3 V20
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3494 0 0
2
45781 4
0
5 4023~
219 681 1348 0 4 22
0 14 15 16 20
0
0 0 624 180
4 4023
-14 -28 14 -20
3 U3B
-8 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 2 3 0
1 U
3507 0 0
2
45781 0
0
7 Pulser~
4 137 1645 0 10 12
0 53 54 55 22 0 0 5 5 6
7
0
0 0 4656 0
0
3 V16
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
5151 0 0
2
45781 10
0
14 Logic Display~
6 766 1607 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3701 0 0
2
45781 9
0
14 Logic Display~
6 577 1627 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8585 0 0
2
45781 8
0
14 Logic Display~
6 415 1633 0 1 2
10 19
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8809 0 0
2
45781 7
0
6 74112~
219 642 1456 0 7 32
0 20 23 15 23 21 16 17
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U8B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 2 8 0
1 U
5993 0 0
2
45781 6
0
6 74112~
219 489 1459 0 7 32
0 20 23 14 23 21 15 18
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U8A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 8 0
1 U
8654 0 0
2
45781 5
0
6 74112~
219 325 1465 0 7 32
0 20 23 22 23 21 14 19
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U7B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 2 7 0
1 U
7223 0 0
2
45781 4
0
7 Pulser~
4 189 1195 0 10 12
0 56 57 58 28 0 0 5 5 6
7
0
0 0 4656 0
0
3 V12
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3641 0 0
2
45781 10
0
14 Logic Display~
6 818 1157 0 1 2
10 25
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3104 0 0
2
45781 9
0
14 Logic Display~
6 629 1177 0 1 2
10 27
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3296 0 0
2
45781 8
0
14 Logic Display~
6 467 1183 0 1 2
10 24
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8534 0 0
2
45781 7
0
6 74112~
219 694 1006 0 7 32
0 30 29 27 29 26 59 25
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U7A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 7 0
1 U
949 0 0
2
45781 6
0
6 74112~
219 541 1009 0 7 32
0 30 29 24 29 26 60 27
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U6B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 6 0
1 U
3371 0 0
2
45781 5
0
6 74112~
219 377 1015 0 7 32
0 30 29 28 29 26 61 24
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U6A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 6 0
1 U
7311 0 0
2
45781 4
0
5 4011~
219 762 904 0 3 22
0 24 25 26
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 5 0
1 U
3409 0 0
2
45781 3
0
5 4011~
219 722 447 0 3 22
0 32 31 33
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 5 0
1 U
3526 0 0
2
45781 0
0
6 74112~
219 337 558 0 7 32
0 37 36 35 36 33 62 34
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U4B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 4 0
1 U
4129 0 0
2
45781 10
0
6 74112~
219 501 552 0 7 32
0 37 36 34 36 33 63 32
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U4A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 4 0
1 U
6278 0 0
2
45781 9
0
6 74112~
219 654 549 0 7 32
0 37 36 32 36 33 64 31
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
3482 0 0
2
45781 8
0
14 Logic Display~
6 427 726 0 1 2
10 34
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8323 0 0
2
45781 7
0
14 Logic Display~
6 589 720 0 1 2
10 32
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3984 0 0
2
45781 6
0
14 Logic Display~
6 778 700 0 1 2
10 31
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7622 0 0
2
45781 5
0
7 Pulser~
4 149 738 0 10 12
0 65 66 67 35 0 0 5 5 6
7
0
0 0 4656 0
0
2 V8
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
816 0 0
2
45781 4
0
5 4023~
219 667 58 0 4 22
0 41 40 39 38
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U3A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 1 3 0
1 U
4656 0 0
2
45781 0
0
7 Pulser~
4 95 349 0 10 12
0 68 69 70 42 0 0 5 5 6
7
0
0 0 4656 0
0
2 V4
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
6356 0 0
2
45781 0
0
14 Logic Display~
6 724 311 0 1 2
10 39
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7479 0 0
2
45781 0
0
14 Logic Display~
6 535 331 0 1 2
10 40
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5690 0 0
2
45781 0
0
14 Logic Display~
6 373 337 0 1 2
10 41
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5617 0 0
2
45781 0
0
6 74112~
219 600 160 0 7 32
0 44 43 40 43 38 71 39
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
3903 0 0
2
45781 0
0
6 74112~
219 447 163 0 7 32
0 44 43 41 43 38 72 40
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
4452 0 0
2
45781 0
0
6 74112~
219 283 169 0 7 32
0 44 43 42 43 38 73 41
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
6282 0 0
2
45781 0
0
108
3 0 2 0 0 8192 0 16 0 0 7 3
849 1723
821 1723
821 1756
6 2 3 0 0 8320 0 18 16 0 0 4
882 1809
915 1809
915 1714
900 1714
0 1 4 0 0 8320 0 0 16 13 0 5
577 1809
577 1743
910 1743
910 1732
900 1732
6 3 5 0 0 4224 0 21 18 0 0 4
707 1806
809 1806
809 1800
822 1800
7 1 6 0 0 8320 0 18 17 0 0 5
876 1791
930 1791
930 2012
943 2012
943 2004
5 0 7 0 0 8320 0 18 0 0 23 3
852 1839
852 1843
677 1844
1 0 2 0 0 8320 0 18 0 0 25 4
852 1764
852 1756
657 1756
657 1753
0 0 8 0 0 8320 0 0 0 9 21 5
817 1791
817 1860
205 1860
205 1817
200 1817
2 4 8 0 0 0 0 18 18 0 0 4
828 1791
814 1791
814 1809
828 1809
7 1 9 0 0 8320 0 21 24 0 0 5
701 1788
788 1788
788 2001
801 2001
801 1993
7 1 10 0 0 8320 0 20 23 0 0 5
548 1791
599 1791
599 2021
612 2021
612 2013
7 1 11 0 0 8320 0 19 22 0 0 5
384 1797
437 1797
437 2027
450 2027
450 2019
6 3 4 0 0 0 0 20 21 0 0 4
554 1809
634 1809
634 1797
647 1797
6 3 12 0 0 4224 0 19 20 0 0 4
390 1815
481 1815
481 1800
494 1800
5 1 7 0 0 0 0 19 1 0 0 5
360 1845
360 1854
216 1854
216 1780
202 1780
3 4 13 0 0 8320 0 19 25 0 0 4
330 1806
210 1806
210 2013
202 2013
0 0 8 0 0 0 0 0 0 18 21 4
644 1806
644 1747
256 1747
256 1803
2 4 8 0 0 0 0 21 21 0 0 4
653 1788
639 1788
639 1806
653 1806
0 0 8 0 0 0 0 0 0 20 21 4
492 1809
492 1750
286 1750
286 1803
2 4 8 0 0 0 0 20 20 0 0 4
500 1791
486 1791
486 1809
500 1809
0 1 8 0 0 0 0 0 2 22 0 4
322 1803
200 1803
200 1837
191 1837
2 4 8 0 0 0 0 19 19 0 0 4
336 1797
322 1797
322 1815
336 1815
0 5 7 0 0 0 0 0 21 24 0 4
510 1849
510 1844
677 1844
677 1836
5 5 7 0 0 0 0 19 20 0 0 4
360 1845
360 1849
524 1849
524 1839
0 1 2 0 0 0 0 0 21 26 0 4
524 1756
524 1753
677 1753
677 1761
1 1 2 0 0 0 0 19 20 0 0 4
360 1770
360 1756
524 1756
524 1764
1 0 14 0 0 12416 0 26 0 0 34 5
705 1357
711 1357
711 1486
359 1486
359 1447
0 2 15 0 0 8320 0 0 26 33 0 5
529 1441
529 1368
720 1368
720 1348
705 1348
6 3 16 0 0 8320 0 31 26 0 0 4
672 1438
715 1438
715 1339
705 1339
7 1 17 0 0 8320 0 31 28 0 0 5
666 1420
753 1420
753 1633
766 1633
766 1625
7 1 18 0 0 8320 0 32 29 0 0 5
513 1423
564 1423
564 1653
577 1653
577 1645
7 1 19 0 0 8320 0 33 30 0 0 5
349 1429
402 1429
402 1659
415 1659
415 1651
6 3 15 0 0 0 0 32 31 0 0 4
519 1441
599 1441
599 1429
612 1429
6 3 14 0 0 0 0 33 32 0 0 4
355 1447
446 1447
446 1432
459 1432
4 0 20 0 0 8192 0 26 0 0 46 3
654 1348
639 1348
639 1385
5 1 21 0 0 8192 0 33 6 0 0 5
325 1477
325 1486
181 1486
181 1412
167 1412
3 4 22 0 0 8320 0 33 27 0 0 4
295 1438
175 1438
175 1645
167 1645
0 0 23 0 0 8320 0 0 0 39 42 4
609 1438
609 1379
221 1379
221 1435
2 4 23 0 0 0 0 31 31 0 0 4
618 1420
604 1420
604 1438
618 1438
0 0 23 0 0 0 0 0 0 41 42 4
457 1441
457 1382
251 1382
251 1435
2 4 23 0 0 0 0 32 32 0 0 4
465 1423
451 1423
451 1441
465 1441
0 1 23 0 0 0 0 0 5 43 0 4
287 1435
165 1435
165 1469
156 1469
2 4 23 0 0 0 0 33 33 0 0 4
301 1429
287 1429
287 1447
301 1447
0 5 21 0 0 8320 0 0 31 45 0 4
475 1481
475 1476
642 1476
642 1468
5 5 21 0 0 0 0 33 32 0 0 4
325 1477
325 1481
489 1481
489 1471
0 1 20 0 0 8192 0 0 31 47 0 4
489 1388
489 1385
642 1385
642 1393
1 1 20 0 0 8320 0 33 32 0 0 4
325 1402
325 1388
489 1388
489 1396
0 1 24 0 0 8320 0 0 41 56 0 3
428 979
428 895
738 895
2 0 25 0 0 8192 0 41 0 0 51 3
738 913
734 913
734 970
3 0 26 0 0 8192 0 41 0 0 63 5
789 904
792 904
792 1023
690 1023
690 1026
7 1 25 0 0 8320 0 38 35 0 0 5
718 970
805 970
805 1183
818 1183
818 1175
0 1 27 0 0 4224 0 0 36 55 0 4
590 973
590 1203
629 1203
629 1195
0 1 24 0 0 0 0 0 37 56 0 4
448 979
448 1209
467 1209
467 1201
3 4 28 0 0 8320 0 40 34 0 0 4
347 988
227 988
227 1195
219 1195
7 3 27 0 0 0 0 39 38 0 0 4
565 973
651 973
651 979
664 979
7 3 24 0 0 0 0 40 39 0 0 4
401 979
498 979
498 982
511 982
0 0 29 0 0 8320 0 0 0 58 61 4
661 988
661 929
273 929
273 985
2 4 29 0 0 0 0 38 38 0 0 4
670 970
656 970
656 988
670 988
0 0 29 0 0 0 0 0 0 60 61 4
509 991
509 932
303 932
303 985
2 4 29 0 0 0 0 39 39 0 0 4
517 973
503 973
503 991
517 991
0 1 29 0 0 0 0 0 8 62 0 4
339 985
217 985
217 1019
208 1019
2 4 29 0 0 0 0 40 40 0 0 4
353 979
339 979
339 997
353 997
0 5 26 0 0 8320 0 0 38 64 0 4
527 1031
527 1026
694 1026
694 1018
5 5 26 0 0 0 0 40 39 0 0 4
377 1027
377 1031
541 1031
541 1021
0 1 30 0 0 4096 0 0 9 67 0 4
377 943
228 943
228 962
219 962
0 1 30 0 0 8192 0 0 38 67 0 4
541 938
541 935
694 935
694 943
1 1 30 0 0 8320 0 40 39 0 0 4
377 952
377 938
541 938
541 946
2 0 31 0 0 8192 0 42 0 0 71 3
698 456
694 456
694 513
0 1 32 0 0 8192 0 0 42 75 0 3
535 516
535 438
698 438
3 0 33 0 0 8192 0 42 0 0 83 5
749 447
752 447
752 566
650 566
650 569
7 1 31 0 0 8320 0 45 48 0 0 5
678 513
765 513
765 726
778 726
778 718
0 1 32 0 0 4224 0 0 47 75 0 4
550 516
550 746
589 746
589 738
0 1 34 0 0 4224 0 0 46 76 0 4
408 522
408 752
427 752
427 744
3 4 35 0 0 8320 0 43 49 0 0 4
307 531
187 531
187 738
179 738
7 3 32 0 0 0 0 44 45 0 0 4
525 516
611 516
611 522
624 522
7 3 34 0 0 0 0 43 44 0 0 4
361 522
458 522
458 525
471 525
0 0 36 0 0 8320 0 0 0 78 81 4
621 531
621 472
233 472
233 528
2 4 36 0 0 0 0 45 45 0 0 4
630 513
616 513
616 531
630 531
0 0 36 0 0 0 0 0 0 80 81 4
469 534
469 475
263 475
263 528
2 4 36 0 0 0 0 44 44 0 0 4
477 516
463 516
463 534
477 534
0 1 36 0 0 0 0 0 11 82 0 4
299 528
177 528
177 562
168 562
2 4 36 0 0 0 0 43 43 0 0 4
313 522
299 522
299 540
313 540
0 5 33 0 0 8320 0 0 45 84 0 4
487 574
487 569
654 569
654 561
5 5 33 0 0 0 0 43 44 0 0 4
337 570
337 574
501 574
501 564
0 1 37 0 0 4096 0 0 10 87 0 4
337 486
188 486
188 505
179 505
0 1 37 0 0 8192 0 0 45 87 0 4
501 481
501 478
654 478
654 486
1 1 37 0 0 8320 0 43 44 0 0 4
337 495
337 481
501 481
501 489
4 0 38 0 0 8192 0 50 0 0 104 5
694 58
698 58
698 177
596 177
596 180
0 3 39 0 0 4096 0 0 50 92 0 5
653 124
653 77
630 77
630 67
643 67
0 2 40 0 0 8192 0 0 50 96 0 3
486 127
486 58
643 58
0 1 41 0 0 8320 0 0 50 97 0 5
313 133
313 190
635 190
635 49
643 49
7 1 39 0 0 8320 0 55 52 0 0 5
624 124
711 124
711 337
724 337
724 329
0 1 40 0 0 4224 0 0 53 96 0 4
496 127
496 357
535 357
535 349
0 1 41 0 0 0 0 0 54 97 0 4
354 133
354 363
373 363
373 355
3 4 42 0 0 8320 0 57 51 0 0 4
253 142
133 142
133 349
125 349
7 3 40 0 0 0 0 56 55 0 0 4
471 127
557 127
557 133
570 133
7 3 41 0 0 0 0 57 56 0 0 4
307 133
404 133
404 136
417 136
0 0 43 0 0 8320 0 0 0 99 102 4
567 142
567 83
179 83
179 139
2 4 43 0 0 0 0 55 55 0 0 4
576 124
562 124
562 142
576 142
0 0 43 0 0 0 0 0 0 101 102 4
415 145
415 86
209 86
209 139
2 4 43 0 0 0 0 56 56 0 0 4
423 127
409 127
409 145
423 145
0 1 43 0 0 0 0 0 14 103 0 4
245 139
123 139
123 173
114 173
2 4 43 0 0 0 0 57 57 0 0 4
259 133
245 133
245 151
259 151
0 5 38 0 0 8320 0 0 55 105 0 4
433 185
433 180
600 180
600 172
5 5 38 0 0 0 0 57 56 0 0 4
283 181
283 185
447 185
447 175
0 1 44 0 0 4096 0 0 15 108 0 4
283 97
134 97
134 116
125 116
0 1 44 0 0 8192 0 0 55 108 0 4
447 92
447 89
600 89
600 97
1 1 44 0 0 8320 0 57 56 0 0 4
283 106
283 92
447 92
447 100
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
118 1689 259 1713
128 1697 248 1713
15 MOD10 asny down
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
83 1322 216 1346
93 1330 205 1346
14 MOD7 asny down
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
135 872 316 896
145 880 305 896
20 MOD 5 Asynchorous up
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
95 415 276 439
105 423 265 439
20 MOD 6 Asynchorous up
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
41 26 222 50
51 34 211 50
20 MOD 7 Asynchorous up
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
