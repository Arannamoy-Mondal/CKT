CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 20 30 100 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
20
13 Logic Switch~
5 141 576 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
45780 0
0
13 Logic Switch~
5 141 496 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
391 0 0
2
45780 0
0
13 Logic Switch~
5 103 218 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3124 0 0
2
45780 0
0
13 Logic Switch~
5 105 158 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3421 0 0
2
45780 0
0
14 Logic Display~
6 608 656 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8157 0 0
2
45780 0
0
14 Logic Display~
6 592 562 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5572 0 0
2
45780 0
0
14 Logic Display~
6 583 487 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8901 0 0
2
45780 0
0
5 4001~
219 479 663 0 3 22
0 3 4 2
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U4A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 4 0
1 U
7361 0 0
2
45780 0
0
5 4001~
219 474 548 0 3 22
0 7 7 6
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U3D
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 3 0
1 U
4747 0 0
2
45780 0
0
5 4001~
219 295 658 0 3 22
0 5 5 4
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U3C
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 3 0
1 U
972 0 0
2
45780 0
0
5 4001~
219 292 579 0 3 22
0 8 5 7
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U3B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 3 0
1 U
3472 0 0
2
45780 0
0
5 4001~
219 289 496 0 3 22
0 8 8 3
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U3A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 3 0
1 U
9998 0 0
2
45780 0
0
5 4011~
219 439 346 0 3 22
0 10 10 9
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 2 0
1 U
3536 0 0
2
45780 0
0
5 4011~
219 431 254 0 3 22
0 15 14 13
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 1 0
1 U
4597 0 0
2
45780 0
0
14 Logic Display~
6 513 334 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3835 0 0
2
45780 0
0
14 Logic Display~
6 506 237 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3670 0 0
2
45780 0
0
14 Logic Display~
6 500 164 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5616 0 0
2
45780 0
0
5 4011~
219 324 341 0 3 22
0 12 11 10
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 1 0
1 U
9323 0 0
2
45780 0
0
5 4011~
219 316 255 0 3 22
0 11 11 14
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 1 0
1 U
317 0 0
2
45780 0
0
5 4011~
219 317 163 0 3 22
0 12 12 15
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 1 0
1 U
3108 0 0
2
45780 0
0
26
3 1 2 0 0 4224 0 8 5 0 0 5
518 663
596 663
596 682
608 682
608 674
0 1 3 0 0 4096 0 0 8 11 0 3
355 496
355 654
466 654
3 2 4 0 0 8336 0 10 8 0 0 5
334 658
334 677
458 677
458 672
466 672
0 2 5 0 0 8192 0 0 10 5 0 3
235 649
235 667
282 667
0 1 5 0 0 8192 0 0 10 9 0 3
177 576
177 649
282 649
3 1 6 0 0 4224 0 9 6 0 0 5
513 548
580 548
580 588
592 588
592 580
0 1 7 0 0 8192 0 0 9 8 0 3
407 579
407 539
461 539
3 2 7 0 0 4224 0 11 9 0 0 4
331 579
453 579
453 557
461 557
1 2 5 0 0 4224 0 1 11 0 0 4
153 576
271 576
271 588
279 588
0 1 8 0 0 8192 0 0 11 13 0 3
189 496
189 570
279 570
3 1 3 0 0 4224 0 12 7 0 0 5
328 496
571 496
571 513
583 513
583 505
0 2 8 0 0 0 0 0 12 13 0 3
250 496
250 505
276 505
1 1 8 0 0 4224 0 2 12 0 0 4
153 496
268 496
268 487
276 487
3 1 9 0 0 4224 0 13 15 0 0 5
466 346
501 346
501 360
513 360
513 352
0 2 10 0 0 8192 0 0 13 16 0 3
385 341
385 355
415 355
3 1 10 0 0 4224 0 18 13 0 0 4
351 341
407 341
407 337
415 337
0 2 11 0 0 8192 0 0 18 23 0 3
148 268
148 350
300 350
0 1 12 0 0 4224 0 0 18 26 0 3
170 158
170 332
300 332
3 1 13 0 0 4224 0 14 16 0 0 5
458 254
494 254
494 263
506 263
506 255
3 2 14 0 0 4224 0 19 14 0 0 4
343 255
399 255
399 263
407 263
0 1 15 0 0 4096 0 0 14 24 0 3
364 163
364 245
407 245
0 1 11 0 0 0 0 0 19 23 0 3
256 268
256 246
292 246
1 2 11 0 0 8320 0 3 19 0 0 5
115 218
115 268
288 268
288 264
292 264
3 1 15 0 0 4224 0 20 17 0 0 5
344 163
488 163
488 190
500 190
500 182
0 2 12 0 0 0 0 0 20 26 0 3
248 158
248 172
293 172
1 1 12 0 0 128 0 4 20 0 0 4
117 158
285 158
285 154
293 154
12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
25 553 54 577
35 561 43 577
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
25 470 54 494
35 478 43 494
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
638 536 691 560
648 544 680 560
4 (OR)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
651 633 712 657
661 641 701 657
5 (And)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
556 329 617 353
566 336 606 352
5 (And)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
627 459 688 483
637 467 677 483
5 (Not)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
18 429 151 473
28 437 140 469
14 3.b)Uni of Nor
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
556 230 609 254
566 238 598 254
4 (OR)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
549 154 610 178
559 162 599 178
5 (Not)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
16 199 45 223
26 207 34 223
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
17 137 46 161
27 145 35 161
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
49 46 190 70
59 54 179 70
15 3.a)Uni Of Nand
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
