CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 1100 2 100 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
24
13 Logic Switch~
5 79 1490 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
45780.6 0
0
13 Logic Switch~
5 70 1406 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
45780.6 0
0
13 Logic Switch~
5 63 669 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
45780.6 0
0
13 Logic Switch~
5 55 591 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3421 0 0
2
45780.6 0
0
13 Logic Switch~
5 98 258 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8157 0 0
2
45780.6 0
0
13 Logic Switch~
5 99 209 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5572 0 0
2
45780.6 0
0
5 4081~
219 644 1328 0 3 22
0 2 3 7
0
0 0 624 180
4 4081
-7 -24 21 -16
3 U5A
-13 -25 8 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
8901 0 0
2
45780.6 0
0
14 Logic Display~
6 1018 1671 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7361 0 0
2
45780.6 0
0
14 Logic Display~
6 727 1678 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4747 0 0
2
45780.6 0
0
14 Logic Display~
6 400 1685 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
972 0 0
2
45780.6 0
0
7 Pulser~
4 96 1650 0 10 12
0 20 21 22 8 0 0 5 5 3
7
0
0 0 4656 0
0
2 V7
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3472 0 0
2
45780.6 0
0
6 74112~
219 800 1458 0 7 32
0 5 6 8 6 5 23 2
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U4A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 4 0
1 U
9998 0 0
2
45780.6 0
0
6 74112~
219 517 1456 0 7 32
0 5 2 8 2 5 24 3
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 3 0
1 U
3536 0 0
2
45780.6 0
0
6 74112~
219 251 1457 0 7 32
0 5 7 8 7 5 25 4
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 3 0
1 U
4597 0 0
2
45780.6 0
0
7 Pulser~
4 149 800 0 10 12
0 26 27 28 14 0 0 5 5 3
7
0
0 0 4656 0
0
2 V6
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3835 0 0
2
45780.6 0
0
14 Logic Display~
6 558 824 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3670 0 0
2
45780.6 0
0
14 Logic Display~
6 327 832 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5616 0 0
2
45780.6 0
0
6 74112~
219 438 646 0 7 32
0 11 12 14 12 11 13 9
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 2 2 0
1 U
9323 0 0
2
45780.6 0
0
6 74112~
219 238 647 0 7 32
0 11 13 14 13 11 29 10
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
317 0 0
2
45780.6 0
0
14 Logic Display~
6 531 374 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3108 0 0
2
45780.6 0
0
14 Logic Display~
6 353 372 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4299 0 0
2
45780.6 0
0
7 Pulser~
4 150 401 0 10 12
0 30 31 32 17 0 0 5 5 3
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
9672 0 0
2
45780.6 0
0
6 74112~
219 473 233 0 7 32
0 18 19 17 19 18 33 15
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
7876 0 0
2
45780.6 0
0
6 74112~
219 264 232 0 7 32
0 18 15 17 15 18 34 16
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
6369 0 0
2
45780.6 0
0
44
0 1 2 0 0 4096 0 0 8 14 0 4
865 1422
865 1697
1018 1697
1018 1689
0 1 3 0 0 4224 0 0 9 17 0 4
582 1420
582 1704
727 1704
727 1696
7 1 4 0 0 8320 0 14 10 0 0 5
275 1421
387 1421
387 1711
400 1711
400 1703
0 1 5 0 0 4224 0 0 12 5 0 3
517 1386
800 1386
800 1395
0 1 5 0 0 0 0 0 13 6 0 4
249 1386
249 1380
517 1380
517 1393
0 1 5 0 0 0 0 0 14 9 0 4
130 1490
130 1386
251 1386
251 1394
0 5 5 0 0 0 0 0 12 8 0 5
517 1472
766 1472
766 1478
800 1478
800 1470
0 5 5 0 0 0 0 0 13 9 0 3
251 1477
517 1477
517 1468
1 5 5 0 0 0 0 1 14 0 0 3
91 1490
251 1490
251 1469
0 4 6 0 0 4112 0 0 12 11 0 4
82 1312
757 1312
757 1440
776 1440
1 2 6 0 0 8320 0 2 12 0 0 5
82 1406
82 1295
762 1295
762 1422
776 1422
4 0 2 0 0 12416 0 13 0 0 14 5
493 1438
444 1438
444 1529
850 1529
850 1422
0 4 7 0 0 4096 0 0 14 15 0 3
222 1328
222 1439
227 1439
2 7 2 0 0 0 0 13 12 0 0 6
493 1420
483 1420
483 1368
875 1368
875 1422
824 1422
3 2 7 0 0 4224 0 7 14 0 0 4
617 1328
213 1328
213 1421
227 1421
7 1 2 0 0 0 0 12 7 0 0 4
824 1422
834 1422
834 1337
662 1337
7 2 3 0 0 0 0 13 7 0 0 4
541 1420
672 1420
672 1319
662 1319
0 3 8 0 0 4224 0 0 12 19 0 4
479 1496
762 1496
762 1431
770 1431
0 3 8 0 0 0 0 0 13 20 0 4
213 1496
479 1496
479 1429
487 1429
4 3 8 0 0 0 0 11 14 0 0 4
126 1650
213 1650
213 1430
221 1430
7 1 9 0 0 8320 0 18 16 0 0 5
462 610
545 610
545 850
558 850
558 842
7 1 10 0 0 8320 0 19 17 0 0 5
262 611
314 611
314 858
327 858
327 850
0 1 11 0 0 4224 0 0 18 24 0 3
238 580
438 580
438 583
0 1 11 0 0 0 0 0 19 27 0 4
176 665
176 576
238 576
238 584
1 0 12 0 0 16512 0 4 0 0 28 6
67 591
67 551
204 551
204 550
381 550
381 612
0 5 11 0 0 0 0 0 18 27 0 3
238 664
438 664
438 658
1 5 11 0 0 0 0 3 19 0 0 4
75 669
75 665
238 665
238 659
2 4 12 0 0 0 0 18 18 0 0 6
414 610
381 610
381 612
378 612
378 628
414 628
6 0 13 0 0 12416 0 18 0 0 30 5
468 628
504 628
504 567
171 567
171 611
2 4 13 0 0 0 0 19 19 0 0 4
214 611
161 611
161 629
214 629
0 3 14 0 0 4224 0 0 18 32 0 4
200 754
401 754
401 619
408 619
4 3 14 0 0 0 0 15 19 0 0 4
179 800
200 800
200 620
208 620
7 1 15 0 0 8192 0 23 20 0 0 5
497 197
518 197
518 400
531 400
531 392
7 1 16 0 0 8320 0 24 21 0 0 5
288 196
340 196
340 398
353 398
353 390
0 3 17 0 0 4224 0 0 23 42 0 4
221 303
425 303
425 206
443 206
0 1 18 0 0 4224 0 0 23 37 0 3
264 137
473 137
473 170
0 1 18 0 0 0 0 0 24 39 0 4
152 258
152 137
264 137
264 169
0 5 18 0 0 0 0 0 23 39 0 3
264 252
473 252
473 245
1 5 18 0 0 0 0 5 24 0 0 3
110 258
264 258
264 244
1 0 19 0 0 16512 0 6 0 0 41 7
111 209
111 119
230 119
230 118
430 118
430 211
435 211
2 4 19 0 0 0 0 23 23 0 0 4
449 197
435 197
435 215
449 215
4 3 17 0 0 0 0 22 24 0 0 4
180 401
221 401
221 205
234 205
4 0 15 0 0 12416 0 24 0 0 44 7
240 214
225 214
225 149
535 149
535 202
502 202
502 197
2 7 15 0 0 0 0 24 23 0 0 6
240 196
230 196
230 164
511 164
511 197
497 197
10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
870 1449 899 1473
880 1457 888 1473
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
597 1456 626 1480
607 1464 615 1480
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
298 1447 327 1471
308 1455 316 1471
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 32
20 1210 297 1234
30 1218 286 1234
32 8.C)Mod 8 Synchronous Up counter
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
491 635 520 659
501 643 509 659
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
265 636 294 660
275 644 283 660
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 34
20 443 313 467
30 451 302 467
34 8.b)Mod 4 Synchronous Down Counter
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
535 227 564 251
545 235 553 251
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
300 229 329 253
310 237 318 253
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 32
5 9 282 33
15 17 271 33
32 8.a)Mod 4 Synchronous Up Counter
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
