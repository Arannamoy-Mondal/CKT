CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 4 100 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
38
13 Logic Switch~
5 188 1637 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7903 0 0
2
45780.2 0
0
13 Logic Switch~
5 188 1757 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7121 0 0
2
45780.2 1
0
13 Logic Switch~
5 191 1842 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4484 0 0
2
45780.2 0
0
13 Logic Switch~
5 205 1126 0 10 11
0 29 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5996 0 0
2
45780.2 1
0
13 Logic Switch~
5 208 1211 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7804 0 0
2
45780.2 0
0
13 Logic Switch~
5 67 310 0 10 11
0 34 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5523 0 0
2
45780.2 0
0
13 Logic Switch~
5 64 225 0 10 11
0 35 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3330 0 0
2
45780.2 0
0
14 Logic Display~
6 1288 2160 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3465 0 0
2
45780.2 0
0
14 Logic Display~
6 995 2170 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8396 0 0
2
45780.2 0
0
14 Logic Display~
6 637 2165 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3685 0 0
2
45780.2 0
0
5 4071~
219 1171 1897 0 3 22
0 6 5 2
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U9C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 9 0
1 U
7849 0 0
2
45780.2 0
0
5 4071~
219 857 1911 0 3 22
0 12 11 3
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U9B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 9 0
1 U
6343 0 0
2
45780.2 0
0
5 4071~
219 547 1905 0 3 22
0 16 15 4
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U9A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 9 0
1 U
7376 0 0
2
45780.2 0
0
5 4081~
219 1063 1944 0 3 22
0 8 7 5
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U8B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 8 0
1 U
9156 0 0
2
45780.2 0
0
5 4081~
219 1053 1861 0 3 22
0 9 10 6
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 8 0
1 U
5776 0 0
2
45780.2 0
0
5 4081~
219 733 1949 0 3 22
0 13 7 11
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U7D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 7 0
1 U
7207 0 0
2
45780.2 0
0
5 4081~
219 729 1880 0 3 22
0 14 10 12
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U7C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 7 0
1 U
4459 0 0
2
45780.2 0
0
5 4081~
219 447 1956 0 3 22
0 17 7 15
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U7B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 7 0
1 U
3760 0 0
2
45780.2 0
0
5 4081~
219 442 1879 0 3 22
0 18 10 16
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 7 0
1 U
754 0 0
2
45780.2 0
0
9 Inverter~
13 280 1631 0 2 22
0 7 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
9767 0 0
2
45780.2 0
0
6 74112~
219 376 1796 0 7 32
0 19 21 20 21 19 17 18
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U5A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 5 0
1 U
7978 0 0
2
45780.2 8
0
6 74112~
219 645 1799 0 7 32
0 19 21 18 21 19 13 14
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U4B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 2 4 0
1 U
3142 0 0
2
45780.2 7
0
6 74112~
219 888 1798 0 7 32
0 19 21 14 21 19 8 9
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U4A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 4 0
1 U
3284 0 0
2
45780.2 6
0
7 Pulser~
4 259 1984 0 10 12
0 36 37 38 20 0 0 5 5 4
8
0
0 0 4656 0
0
2 V9
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
659 0 0
2
45780.2 5
0
6 74112~
219 393 1165 0 7 32
0 28 29 27 29 28 24 26
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 2 3 0
1 U
3800 0 0
2
45780.2 8
0
6 74112~
219 662 1168 0 7 32
0 28 29 26 29 28 23 25
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 3 0
1 U
6792 0 0
2
45780.2 7
0
6 74112~
219 905 1167 0 7 32
0 28 29 25 29 28 22 39
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
3701 0 0
2
45780.2 6
0
7 Pulser~
4 276 1353 0 10 12
0 40 41 42 27 0 0 5 5 4
8
0
0 0 4656 0
0
2 V6
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
6316 0 0
2
45780.2 5
0
14 Logic Display~
6 491 991 0 1 2
10 24
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8734 0 0
2
45780.2 4
0
14 Logic Display~
6 725 995 0 1 2
10 23
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7988 0 0
2
45780.2 3
0
14 Logic Display~
6 1000 989 0 1 2
10 22
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3217 0 0
2
45780.2 2
0
14 Logic Display~
6 859 88 0 1 2
10 30
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3965 0 0
2
45780.2 0
0
14 Logic Display~
6 584 94 0 1 2
10 31
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8239 0 0
2
45780.2 0
0
14 Logic Display~
6 350 90 0 1 2
10 32
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
828 0 0
2
45780.2 0
0
7 Pulser~
4 135 452 0 10 12
0 43 44 45 33 0 0 5 5 4
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
6187 0 0
2
45780.2 0
0
6 74112~
219 764 266 0 7 32
0 34 35 31 35 34 46 30
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
7107 0 0
2
45780.2 0
0
6 74112~
219 521 267 0 7 32
0 34 35 32 35 34 47 31
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
6433 0 0
2
45780.2 0
0
6 74112~
219 252 264 0 7 32
0 34 35 33 35 34 48 32
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
8559 0 0
2
45780.2 0
0
73
3 1 2 0 0 8320 0 11 8 0 0 5
1204 1897
1275 1897
1275 2186
1288 2186
1288 2178
3 1 3 0 0 8320 0 12 9 0 0 5
890 1911
982 1911
982 2196
995 2196
995 2188
3 1 4 0 0 8320 0 13 10 0 0 5
580 1905
624 1905
624 2191
637 2191
637 2183
3 2 5 0 0 4224 0 14 11 0 0 4
1084 1944
1150 1944
1150 1906
1158 1906
3 1 6 0 0 4224 0 15 11 0 0 4
1074 1861
1150 1861
1150 1888
1158 1888
0 2 7 0 0 8336 0 0 14 37 0 5
201 1637
201 2121
1031 2121
1031 1953
1039 1953
6 1 8 0 0 8320 0 23 14 0 0 4
918 1780
1024 1780
1024 1935
1039 1935
7 1 9 0 0 4224 0 23 15 0 0 4
912 1762
1016 1762
1016 1852
1029 1852
0 2 10 0 0 4224 0 0 15 15 0 4
697 1666
1021 1666
1021 1870
1029 1870
3 2 11 0 0 4224 0 16 12 0 0 4
754 1949
836 1949
836 1920
844 1920
3 1 12 0 0 4224 0 17 12 0 0 4
750 1880
836 1880
836 1902
844 1902
6 1 13 0 0 8320 0 22 16 0 0 4
675 1781
701 1781
701 1940
709 1940
0 2 7 0 0 0 0 0 16 37 0 7
200 1637
200 2069
419 2069
419 2013
701 2013
701 1958
709 1958
0 1 14 0 0 4096 0 0 17 28 0 3
685 1763
685 1871
705 1871
0 2 10 0 0 0 0 0 17 20 0 4
403 1644
697 1644
697 1889
705 1889
3 2 15 0 0 4224 0 18 13 0 0 4
468 1956
526 1956
526 1914
534 1914
3 1 16 0 0 4224 0 19 13 0 0 4
463 1879
526 1879
526 1896
534 1896
0 2 7 0 0 0 0 0 18 37 0 5
215 1637
215 2029
415 2029
415 1965
423 1965
6 1 17 0 0 8320 0 21 18 0 0 4
406 1778
411 1778
411 1947
423 1947
2 2 10 0 0 0 0 20 19 0 0 4
301 1631
403 1631
403 1888
418 1888
0 1 18 0 0 4096 0 0 19 29 0 3
420 1760
420 1870
418 1870
0 1 19 0 0 4096 0 0 23 23 0 3
645 1723
888 1723
888 1735
0 1 19 0 0 8320 0 0 22 24 0 4
311 1725
311 1718
645 1718
645 1736
0 1 19 0 0 0 0 0 21 27 0 4
251 1842
251 1725
376 1725
376 1733
0 5 19 0 0 0 0 0 23 26 0 3
645 1826
888 1826
888 1810
0 5 19 0 0 0 0 0 22 27 0 3
376 1831
645 1831
645 1811
1 5 19 0 0 0 0 3 21 0 0 3
203 1842
376 1842
376 1808
7 3 14 0 0 4224 0 22 23 0 0 4
669 1763
850 1763
850 1771
858 1771
7 3 18 0 0 4224 0 21 22 0 0 4
400 1760
602 1760
602 1772
615 1772
4 3 20 0 0 8320 0 24 21 0 0 4
289 1984
338 1984
338 1769
346 1769
0 4 21 0 0 12288 0 0 23 32 0 6
607 1803
611 1803
611 1816
850 1816
850 1780
864 1780
0 4 21 0 0 8192 0 0 22 33 0 5
343 1778
343 1812
607 1812
607 1781
621 1781
0 4 21 0 0 0 0 0 21 36 0 3
301 1757
301 1778
352 1778
0 2 21 0 0 0 0 0 23 35 0 5
607 1728
607 1731
850 1731
850 1762
864 1762
0 2 21 0 0 8320 0 0 22 36 0 5
342 1757
342 1728
607 1728
607 1763
621 1763
1 2 21 0 0 0 0 2 21 0 0 4
200 1757
338 1757
338 1760
352 1760
1 1 7 0 0 0 0 1 20 0 0 4
200 1637
257 1637
257 1631
265 1631
6 1 22 0 0 8320 0 27 31 0 0 3
935 1149
1000 1149
1000 1007
6 1 23 0 0 8320 0 26 30 0 0 3
692 1150
725 1150
725 1013
6 1 24 0 0 8320 0 25 29 0 0 3
423 1147
491 1147
491 1009
7 3 25 0 0 4224 0 26 27 0 0 4
686 1132
867 1132
867 1140
875 1140
7 3 26 0 0 4224 0 25 26 0 0 4
417 1129
619 1129
619 1141
632 1141
4 3 27 0 0 8320 0 28 25 0 0 4
306 1353
355 1353
355 1138
363 1138
0 1 28 0 0 8192 0 0 27 45 0 4
662 1092
662 1096
905 1096
905 1104
0 1 28 0 0 8320 0 0 26 46 0 4
393 1080
393 1092
662 1092
662 1105
0 1 28 0 0 0 0 0 25 52 0 4
268 1213
268 1080
393 1080
393 1102
0 4 29 0 0 12288 0 0 27 48 0 6
624 1165
628 1165
628 1176
867 1176
867 1149
881 1149
0 4 29 0 0 8320 0 0 26 49 0 5
340 1147
340 1182
624 1182
624 1150
638 1150
0 4 29 0 0 0 0 0 25 55 0 3
302 1126
302 1147
369 1147
0 5 28 0 0 0 0 0 27 51 0 3
662 1187
905 1187
905 1179
0 5 28 0 0 0 0 0 26 52 0 3
393 1196
662 1196
662 1180
1 5 28 0 0 0 0 5 25 0 0 4
220 1211
220 1213
393 1213
393 1177
0 2 29 0 0 0 0 0 27 54 0 4
624 1101
867 1101
867 1131
881 1131
0 2 29 0 0 0 0 0 26 55 0 5
359 1126
359 1097
624 1097
624 1132
638 1132
1 2 29 0 0 0 0 4 25 0 0 4
217 1126
355 1126
355 1129
369 1129
7 1 30 0 0 8320 0 36 32 0 0 3
788 230
859 230
859 106
0 1 31 0 0 4096 0 0 33 59 0 2
584 231
584 112
0 1 32 0 0 4096 0 0 34 60 0 2
350 228
350 108
7 3 31 0 0 4224 0 37 36 0 0 4
545 231
726 231
726 239
734 239
7 3 32 0 0 4224 0 38 37 0 0 4
276 228
478 228
478 240
491 240
4 3 33 0 0 8320 0 35 38 0 0 4
165 452
214 452
214 237
222 237
0 1 34 0 0 8192 0 0 36 63 0 4
521 191
521 195
764 195
764 203
0 1 34 0 0 8320 0 0 37 64 0 4
252 179
252 191
521 191
521 204
0 1 34 0 0 0 0 0 38 70 0 4
127 312
127 179
252 179
252 201
0 4 35 0 0 12288 0 0 36 66 0 6
483 264
487 264
487 275
726 275
726 248
740 248
0 4 35 0 0 8320 0 0 37 67 0 5
199 246
199 281
483 281
483 249
497 249
0 4 35 0 0 0 0 0 38 73 0 3
161 225
161 246
228 246
0 5 34 0 0 0 0 0 36 69 0 3
521 286
764 286
764 278
0 5 34 0 0 0 0 0 37 70 0 3
252 295
521 295
521 279
1 5 34 0 0 0 0 6 38 0 0 4
79 310
79 312
252 312
252 276
0 2 35 0 0 0 0 0 36 72 0 4
483 200
726 200
726 230
740 230
0 2 35 0 0 0 0 0 37 73 0 5
218 225
218 196
483 196
483 231
497 231
1 2 35 0 0 0 0 7 38 0 0 4
76 225
214 225
214 228
228 228
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 32
76 1532 353 1556
86 1540 342 1556
32 7.C)Asynchronous UP-Down Counter
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 33
18 6 303 30
28 14 292 30
33 7.a)Mod 8 asynchronous Up Counter
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 35
47 845 348 869
57 853 337 869
35 7.b)Mod 8 asynchronous Down Counter
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
