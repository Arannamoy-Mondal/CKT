CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
13
13 Logic Switch~
5 109 527 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8748 0 0
2
45780.1 0
0
13 Logic Switch~
5 112 471 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7168 0 0
2
45780.1 0
0
13 Logic Switch~
5 75 263 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
631 0 0
2
45780.1 0
0
13 Logic Switch~
5 70 217 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9466 0 0
2
45780.1 0
0
13 Logic Switch~
5 68 163 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3266 0 0
2
45780.1 0
0
14 Logic Display~
6 477 545 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7693 0 0
2
45780.1 0
0
14 Logic Display~
6 476 476 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3723 0 0
2
45780.1 0
0
7 Pulser~
4 106 621 0 10 12
0 13 14 4 15 0 0 5 5 4
8
0
0 0 4656 0
0
2 V5
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3440 0 0
2
45780.1 0
0
6 74LS74
17 273 500 0 12 25
0 4 6 5 5 16 17 18 19 3
2 20 21
0
0 0 4848 0
6 74LS74
-21 -60 21 -52
2 U2
-7 -61 7 -53
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 3 2 4 1 11 12 10 13 5
6 9 8 3 2 4 1 11 12 10
13 5 6 9 8 0
65 0 0 512 0 0 0 0
1 U
6263 0 0
2
45780.1 0
0
7 Pulser~
4 130 348 0 10 12
0 22 23 24 7 0 0 5 5 4
8
0
0 0 4656 0
0
2 V4
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
4900 0 0
2
45780.1 0
0
14 Logic Display~
6 398 215 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8783 0 0
2
45780.1 0
0
14 Logic Display~
6 395 151 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3221 0 0
2
45780.1 0
0
6 74LS76
104 221 187 0 14 29
0 12 11 7 10 10 25 26 27 28
29 9 8 30 31
0
0 0 4848 0
6 74LS76
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=13;
130 %D [%5bi %13bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 16 1 2 3 9 12 6 7
8 15 14 11 10 4 16 1 2 3
9 12 6 7 8 15 14 11 10 0
65 0 0 512 0 0 0 0
1 U
3215 0 0
2
45780.1 0
0
13
10 1 2 0 0 4224 0 9 6 0 0 5
311 482
459 482
459 571
477 571
477 563
9 1 3 0 0 4224 0 9 7 0 0 5
305 473
464 473
464 502
476 502
476 494
3 1 4 0 0 8320 0 8 9 0 0 4
130 612
222 612
222 464
241 464
0 3 5 0 0 8192 0 0 9 5 0 3
179 527
179 482
235 482
1 4 5 0 0 4224 0 1 9 0 0 4
121 527
227 527
227 491
235 491
1 2 6 0 0 4224 0 2 9 0 0 4
124 471
227 471
227 473
241 473
4 3 7 0 0 8320 0 10 13 0 0 4
160 348
165 348
165 169
183 169
12 1 8 0 0 4224 0 13 11 0 0 5
259 160
378 160
378 241
398 241
398 233
11 1 9 0 0 4224 0 13 12 0 0 5
253 151
383 151
383 177
395 177
395 169
0 4 10 0 0 4096 0 0 13 11 0 3
118 263
118 178
183 178
1 5 10 0 0 4224 0 3 13 0 0 4
87 263
175 263
175 187
183 187
1 2 11 0 0 4224 0 4 13 0 0 4
82 217
170 217
170 160
189 160
1 1 12 0 0 8336 0 5 13 0 0 5
80 163
80 150
175 150
175 151
189 151
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
21 397 210 421
31 405 199 421
21 6.c)D Flip-flop(7474)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 24
25 29 238 53
35 37 227 53
24 6.a)b)Jk Flip-Flop(7476)
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
