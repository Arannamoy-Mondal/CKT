CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 136 241 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
45779.9 0
0
13 Logic Switch~
5 138 171 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
45779.9 0
0
5 4001~
219 228 637 0 3 22
0 4 3 2
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U6A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 6 0
1 U
3124 0 0
2
45779.9 0
0
5 4011~
219 383 567 0 3 22
0 4 3 5
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 5 0
1 U
3421 0 0
2
45779.9 0
0
14 Logic Display~
6 629 647 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8157 0 0
2
45779.9 0
0
5 4030~
219 242 503 0 3 22
0 4 3 6
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U4A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
5572 0 0
2
45779.9 0
0
14 Logic Display~
6 623 566 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8901 0 0
2
45779.9 0
0
14 Logic Display~
6 616 489 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7361 0 0
2
45779.9 0
0
14 Logic Display~
6 611 404 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4747 0 0
2
45779.9 0
0
9 Inverter~
13 281 399 0 2 22
0 4 7
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
972 0 0
2
45779.9 0
0
5 4071~
219 355 321 0 3 22
0 4 3 8
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
3472 0 0
2
45779.9 0
0
14 Logic Display~
6 597 277 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9998 0 0
2
45779.9 0
0
14 Logic Display~
6 590 181 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3536 0 0
2
45779.9 0
0
5 4081~
219 345 187 0 3 22
0 4 3 9
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
4597 0 0
2
45779.9 0
0
17
3 1 2 0 0 4224 0 3 5 0 0 5
267 637
617 637
617 673
629 673
629 665
0 2 3 0 0 4224 0 0 3 16 0 3
207 241
207 646
215 646
0 1 4 0 0 4224 0 0 3 17 0 3
168 171
168 628
215 628
3 1 5 0 0 4224 0 4 7 0 0 5
410 567
611 567
611 592
623 592
623 584
0 2 3 0 0 0 0 0 4 16 0 6
246 241
246 440
306 440
306 575
359 575
359 576
0 1 4 0 0 16 0 0 4 17 0 5
306 171
306 428
354 428
354 558
359 558
3 1 6 0 0 4224 0 6 8 0 0 5
275 503
604 503
604 515
616 515
616 507
0 2 3 0 0 128 0 0 6 16 0 5
151 241
151 231
151 231
151 512
226 512
0 1 4 0 0 128 0 0 6 17 0 3
184 171
184 494
226 494
2 1 7 0 0 4224 0 10 9 0 0 5
302 399
599 399
599 430
611 430
611 422
0 1 4 0 0 128 0 0 10 17 0 3
227 171
227 399
266 399
3 1 8 0 0 4224 0 11 12 0 0 3
388 321
597 321
597 295
0 2 3 0 0 128 0 0 11 16 0 3
173 241
173 330
342 330
0 1 4 0 0 0 0 0 11 17 0 3
197 171
197 312
342 312
3 1 9 0 0 4224 0 14 13 0 0 5
366 187
578 187
578 207
590 207
590 199
1 2 3 0 0 128 0 1 14 0 0 4
148 241
313 241
313 196
321 196
1 1 4 0 0 128 0 2 14 0 0 4
150 171
313 171
313 178
321 178
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
86 217 111 241
94 225 102 241
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
88 153 117 177
98 161 106 177
1 A
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
